module primeiro_codigo (
	output [7:0] LED
);

assign LED = 8'h55;

endmodule
